module hello_world_example;

initial begin
  $display("Hello, World!");
end

endmodule
